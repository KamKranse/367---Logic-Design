library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CPU is
  port(clock    : in  std_logic;
       reset    : in  std_logic;
       from_mem : in  std_logic_vector(7 downto 0);
       write    : out std_logic;
       to_mem   : out std_logic_vector(7 downto 0);
       address  : out std_logic_vector(7 downto 0));
  end entity;
  
  
  architecture CPU_arch of CPU is 
  
  component data_path is
  port(clock       : in  std_logic;
       reset       : in  std_logic;
       IR_Load     : in  std_logic;
       MAR_Load    : in  std_logic;
       PC_Load     : in  std_logic;
       PC_Inc      : in  std_logic;
       A_Load      : in  std_logic;
       B_Load      : in  std_logic;
       ALU_Sel     : in  std_logic_vector(2 downto 0);
       CCR_Load    : in  std_logic;
       Bus2_Sel    : in  std_logic_vector(1 downto 0);
       Bus1_Sel    : in  std_logic_vector(1 downto 0);
       from_memory : in  std_logic_vector(7 downto 0);
       CCR_Result  : out std_logic_vector(3 downto 0);
       IR          : out std_logic_vector(7 downto 0);
       address     : out std_logic_vector(7 downto 0);
       to_memory   : out std_logic_vector(7 downto 0));
  end component;

  component control_unit is
	port	(Clock       : in  std_logic;
	      Reset       : in  std_logic;
	      CCR_Results : in  std_logic_vector(3 downto 0);
	      IR          : in  std_logic_vector(7 downto 0);
	      IR_Load     : out std_logic;
	      MAR_Load    : out std_logic;
	      PC_Load     : out std_logic;
	      PC_Inc      : out std_logic;
	      A_Load      : out std_logic;
	      B_Load      : out std_logic;
	      ALU_Sel     : out std_logic_vector(2 downto 0);
	      CCR_Load    : out std_logic;
	      Bus1_Sel    : out std_logic_vector(1 downto 0);
	      Bus2_Sel    : out std_logic_vector(1 downto 0);
	      write       : out std_logic);
  end component;
  
  signal  IR_Load, MAR_Load, PC_Load, PC_Inc, A_Load, B_Load, CCR_Load  : std_logic;
  signal  ALU_Sel                                                       : std_logic_vector(2 downto 0);
  signal  bus1_sel, bus2_sel                                            : std_logic_vector(1 downto 0);
  signal  IR                                                            : std_logic_vector(7 downto 0);
  signal  CCR_result                                                    : std_logic_vector(3 downto 0);
    
  
  begin

    CU  : control_unit port map(clock, reset, CCR_Result, IR,       IR_Load, MAR_Load, PC_Load, PC_Inc, A_Load,  B_Load,   ALU_Sel,  CCR_Load, bus1_sel, bus2_sel,   write);
    
    DP  : data_path port map   (clock, reset, IR_Load,    MAR_Load, PC_Load, PC_Inc,   A_Load,  B_Load, ALU_Sel, CCR_Load, bus2_sel, bus1_sel, from_mem, CCR_Result, IR, address, to_mem);
  
  end architecture;
  
     
       
       
